`ifndef SIGN_EXTENDER_TYPES
`define SIGN_EXTENDER_TYPES

typedef enum logic {
  TYPE_I = 1'b0,
  ERROR = 1'b1
} sign_extender_control_t;

`endif // SIGN_EXTENDER_TYPES